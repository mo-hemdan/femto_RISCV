`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/23/2020 02:12:37 PM
// Design Name: 
// Module Name: inst_mem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module InstMem (input [6:0] addr, output [31:0] data_out);
 reg [31:0] mem [0:127];
 assign data_out = mem[addr];
 initial begin
 /*mem[3:0] = 32'h004e80b7;
 mem[1] = 32'h00000033;
 mem[2] = 32'h00000033;
 mem[3] = 32'h00000033;
 mem[4] = 32'h0300e093;
 mem[5] = 32'h00000033;
 mem[6] = 32'h00000033;
 mem[7] = 32'h00000033;
 mem[8] = 32'h01efe117;
 mem[9] = 32'h00000033;
 mem[10] = 32'h00000033;
 mem[11] = 32'h00000033;
 mem[12] = 32'h00000183;
 mem[13] = 32'h00000033;
 mem[14] = 32'h00000033;
 mem[15] = 32'h00000033;
 mem[16] = 32'h00001203;
 mem[17] = 32'h00000033;
 mem[18] = 32'h00000033;
 mem[19] = 32'h00000033;
 mem[20] = 32'h00002283;
 mem[21] = 32'h00000033;
 mem[22] = 32'h00000033;
 mem[23] = 32'h00000033;
 mem[24] = 32'h00500223;
 mem[25] = 32'h00000033;
 mem[26] = 32'h00000033;
 mem[27] = 32'h00000033;
 mem[28] = 32'h00501423;
 mem[29] = 32'h00000033;
 mem[30] = 32'h00000033;
 mem[31] = 32'h00000033;
 mem[32] = 32'h00502623;
 mem[33] = 32'h00000033;
 mem[34] = 32'h00000033;
 mem[35] = 32'h00000033;
 mem[36] = 32'h00008133;
 mem[37] = 32'h00000033;
 mem[38] = 32'h00000033;
 mem[39] = 32'h00000033;
 mem[40] = 32'h40110133;
 mem[41] = 32'h00000033;
 mem[42] = 32'h00000033;
 mem[43] = 32'h00000033;
 mem[44] = 32'h00329333;
 mem[45] = 32'h00000033;
 mem[46] = 32'h00000033;
 mem[47] = 32'h00000033;
 mem[48] = 32'h0032d3b3;
 mem[49] = 32'h00000033;
 mem[50] = 32'h00000033;
 mem[51] = 32'h00000033;
 mem[52] = 32'hf3800393;
 mem[53] = 32'h00000033;
 mem[54] = 32'h00000033;
 mem[55] = 32'h00000033;
 mem[56] = 32'h4033d3b3;
 mem[57] = 32'h00000033;
 mem[58] = 32'h00000033;
 mem[59] = 32'h00000033;
 mem[60] = 32'h00712433;
 mem[61] = 32'h00000033;
 mem[62] = 32'h00000033;
 mem[63] = 32'h00000033;
 mem[64] = 32'h007334b3;
 mem[65] = 32'h00000033;
 mem[66] = 32'h00000033;
 mem[67] = 32'h00000033;
 mem[68] = 32'h006344b3;
 mem[69] = 32'h00000033;
 mem[70] = 32'h00000033;
 mem[71] = 32'h00000033;
 mem[72] = 32'hfff00313;
 mem[73] = 32'h00000033;
 mem[74] = 32'h00000033;
 mem[75] = 32'h00000033;
 mem[76] = 32'h0060e4b3;
 mem[77] = 32'h00000033;
 mem[78] = 32'h00000033;
 mem[79] = 32'h00000033;
 mem[80] = 32'h0000f0b3;
 mem[81] = 32'h00000033;
 mem[82] = 32'h00000033;
 mem[83] = 32'h00000033;*/
/*
   mem[0] = 32'h004e80b7;
   mem[1]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[2]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[3]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[4] = 32'h00000033;
   mem[5]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[6]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[7]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[8] = 32'h00000033;
   mem[9]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[10]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[11]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[12] = 32'h00000033;
   mem[13]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[14]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[15]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[16] = 32'h0300e093;
   mem[17]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[18]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[19]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[20] = 32'h00000033;
   mem[21]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[22]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[23]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[24] = 32'h00000033;
   mem[25]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[26]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[27]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[28] = 32'h00000033;
   mem[29]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[30]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[31]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[32] = 32'h01efe117;
   mem[33]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[34]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[35]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[36] = 32'h00000033;
   mem[37]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[38]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[39]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[40] = 32'h00000033;
   mem[41]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[42]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[43]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[44] = 32'h00000033;
   mem[45] =32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[46] = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[47]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[48] = 32'h00000183;
   mem[49]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[50]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[51]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[52] = 32'h00000033;
   mem[53]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[54]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[55]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[56] = 32'h00000033;
   mem[57]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[58]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[59]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[60] = 32'h00000033;
   mem[61]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[62]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[63]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[64] = 32'h00001203;
   mem[65]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[66]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[67]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[68] = 32'h00000033;
   mem[69]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[70]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[71]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[72] = 32'h00000033;
   mem[73]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[74]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[75]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[76] = 32'h00000033;
   mem[77]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[78]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[79]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[80] = 32'h00002283;
   mem[81]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[82]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[83]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[84] = 32'h00000033;
   mem[85]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[86]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[87]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[88] = 32'h00000033;
   mem[89]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[90]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[91]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[92] = 32'h00000033;
   mem[93]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[94]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[95]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[96] = 32'h00500223;
   mem[97]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[98]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[99]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[100] = 32'h00000033;
   mem[101]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[102]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[103]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[104] = 32'h00000033;
   mem[105]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[106]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[107]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[108] = 32'h00000033;
   mem[109]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[110]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[111]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[112] = 32'h00501423;
   mem[113]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[114]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[115]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[116] = 32'h00000033;
   mem[117]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[118]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[119]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[120]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[121] = 32'h00000033;
   mem[122]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[123]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[124]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[125] = 32'h00000033;
   mem[126]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[127]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[128]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[129] = 32'h00502623;
   mem[130]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[131]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[132]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[133] = 32'h00000033;
   mem[134]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[135]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[136]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[137] = 32'h00000033;
   mem[138]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[139]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[140]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[141]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[142] = 32'h00000033;
   mem[143]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[144]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[145]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[146] = 32'h00008133;
   mem[147]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[148]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[149]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[150] = 32'h00000033;
   mem[151]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[152]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[153]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[154] = 32'h00000033;
   mem[155]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[156]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[157]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[158] = 32'h00000033;
   mem[159]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[160]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[161]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[162] = 32'h40110133;
   mem[163]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[164]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[165]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[166]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[167] = 32'h00000033;
   mem[168]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[169]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[170]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[171] = 32'h00000033;
   mem[172]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[173]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[174]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[175] = 32'h00000033;
   mem[176]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[177]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[178]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[179] = 32'h00329333;
   mem[180]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[181]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[182]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[183] = 32'h00000033;
   mem[184]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[185]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[186]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[187] = 32'h00000033;
   mem[188]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[189]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[190]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[191]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[192] = 32'h00000033;
   mem[193]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[194]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0  //mem[195]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[195] = 32'h0032d3b3;
   mem[196]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[197]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0  //mem[199]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[198] = 32'h00000033;
   mem[199]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[200]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[201]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[202] = 32'h00000033;
   mem[203]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[204]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[205]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[206] = 32'h00000033;
   mem[207]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[208]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[209]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[210] = 32'hf3800393;
   mem[211]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[212]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[213]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[214] = 32'h00000033;
   mem[215]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[216]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[217]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[218] = 32'h00000033;
   mem[219]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[220]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[221]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[222] = 32'h00000033;
   mem[223]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[224]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[225]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[226] = 32'h4033d3b3;
   mem[227]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[228]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[229]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[230] = 32'h00000033;
   mem[2]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[230]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[231]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[232] = 32'h00000033;
   mem[233]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[234]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[235]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[236] = 32'h00000033;
   mem[237]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[238]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[239]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[240] = 32'h00712433;
   mem[241]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[242]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[243]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[244] = 32'h00000033;
   mem[245]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[246]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[247]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[248] = 32'h00000033;
   mem[249]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[250]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[251]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[252] = 32'h00000033;
   mem[253]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[254]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[255]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[256] = 32'h007334b3;
   mem[257]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[258]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[259]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[260] = 32'h00000033;
   mem[261]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[262]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[263]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[264] = 32'h00000033;
   mem[265]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[266]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[267]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[268] = 32'h00000033;
   mem[269]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[270]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[271]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[272] = 32'h006344b3;
   mem[273]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[274]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[275]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[276] = 32'h00000033;
   mem[277]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[278]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[279]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[280] = 32'h00000033;
   mem[281]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[282]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[283]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[284] = 32'h00000033;
   mem[285]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[286]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[287]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[288] = 32'hfff00313;
   mem[289]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[290]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[291]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[292] = 32'h00000033;
   mem[293]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[294]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[295]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[296]= 32'h00000033;
   mem[297]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[298]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[299]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[300] = 32'h00000033;
   mem[301]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[302]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[303]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[304] = 32'h0060e4b3;
   mem[305]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[306]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[307]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[308] = 32'h00000033;
   mem[309]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[310]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[311]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[312] = 32'h00000033;
   mem[313]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[314]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[315]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[316] = 32'h00000033;
   mem[317]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[318]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[319]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[320] = 32'h0000f0b3;
   mem[321]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[322]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[323]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[324] = 32'h00000033;
   mem[325]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[326]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[327]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[328] = 32'h00000033;
   mem[329]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[330]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[331]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[332] = 32'h00000033;
   mem[333]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[334]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
   mem[335]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0*/
  /*mem[0]=32'b00000000000000000000000010110011;
  mem[1]=32'b00000000110100000000000010010011;
  mem[2]=32'b00000000010100001110000010010011;
  mem[3]=32'b00000000010100001100000100010011;
  mem[4]=32'b11111111011100010000000100010011;
  mem[5]=32'b00000000011000010010000110010011;
  mem[6]=32'b00000000100100010010001000010011;
  mem[7]=32'b00000000011000010011001100010011;
  mem[8]=32'b00000000001000010001001110010011;
  mem[9]=32'b00000000001000010101010000010011;
  mem[10]=32'b01000000001000010101010010010011;
 */
 

// i don't know what program is this 

  //mem[0]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
  //mem[1]=32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0)
  //mem[2]=32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0)
  //mem[3]=32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0)
  //mem[4]=32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2
  //mem[5]=32'b0_000000_00011_00100_000_0100_0_1100011 ; //beq x4, x3, 4
  //mem[6]=32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2
  //mem[7]=32'b0000000_00010_00011_000_00101_0110011 ; //add x5, x3, x2
  //mem[8]=32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0)
  //mem[9]=32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)
  //mem[10]=32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1
  //mem[11]=32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2
  //mem[12]=32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2
  //mem[13]=32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1
 end
 
endmodule
